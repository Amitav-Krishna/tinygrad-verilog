module tb_layer;
  reg clk;
  reg start;

  reg signed [31:0] x_vals;
  reg signed [63:0] w_vals;
  reg signed [31:0] b_vals;

  wire signed [31:0] y;
  wire done;

  layer #(
    .N(2),
    .M(2)
   ) uut (
    .clk(clk),
    .start(start),
    .x(x_vals),
    .w(w_vals),
    .b(b_vals),
    .y(y),
    .done(done)
  );

  always #5 clk = ~clk;

  // ~ is the not operator, which makes clock flip every 5 time units.
  
  // Helper functions
  function real q8_to_real;
      input signed [15:0] q;
      begin
          q8_to_real = $itor(q) / 256.0;
      end
  endfunction

  function signed [15:0] real_to_q8;
      input real r;
      begin
          real_to_q8 = $rtoi(r * 256.0);
      end
  endfunction

  initial begin
    $display("=== Layer Unit Test ===");

     // Initialize vectors (Q8.8 fixed point)
     x_vals = {
	       real_to_q8(2.0),
	       real_to_q8(1.0)
	       };

    
     w_vals = {
	       real_to_q8(0.4), real_to_q8(0.3),

	       real_to_q8(0.7), real_to_q8(0.5)
	       };

    // Zero biases
    b_vals = {
      real_to_q8(1.2),
      real_to_q8(0.7)
    };

    clk = 0;
    start = 0;

    #20;
    start = 1;
    #10;
    start = 0;

     #200;

     $display("Inputs:  [%.3f, %.3f]",
	      q8_to_real(x_vals[15:0]),
	      q8_to_real(x_vals[31:16])
	      );
     

     $display("Outputs: [%.3f, %.3f]",
	      q8_to_real(y[15:0]),
	      q8_to_real(y[31:16])
	      );
     


     $display("Done: %b", done);

  end
endmodule

